/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */
`default_nettype none

module tt_um_uwasic_onboarding_Hugh_Ding (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  // assign uo_out  = 8'b11111111;  // Example: ou_out is the sum of ui_in and uio_in 
  // assign uio_out = 0;
  
  assign uio_oe  = 8'hFF;

  wire [7:0] en_reg_out_7_0;
  wire [7:0] en_reg_out_15_8;
  wire [7:0] en_reg_pwm_7_0;
  wire [7:0] en_reg_pwm_15_8;
  wire [7:0] pwm_duty_cycle;

  spi_peripheral spi_peripheral_inst (
    .SCLK(ui_in[0]),
    .nCS(ui_in[2]),
    .COPI(ui_in[1]),
    .clk(clk),
    .rst_n(rst_n),
    .EN_REG_OUT_7_0(en_reg_out_7_0),
    .EN_REG_OUT_15_8(en_reg_out_15_8),
    .EN_REG_PWM_7_0(en_reg_pwm_7_0),
    .EN_REG_PWM_15_8(en_reg_pwm_15_8),
    .PWM_DUTY_CYCLE(pwm_duty_cycle)
  );

   pwm_peripheral pwm_peripheral_inst (
    .clk(clk),
    .rst_n(rst_n),
    .en_reg_out_7_0(en_reg_out_7_0),
    .en_reg_out_15_8(en_reg_out_15_8),
    .en_reg_pwm_7_0(en_reg_pwm_7_0),
    .en_reg_pwm_15_8(en_reg_pwm_15_8),
    .pwm_duty_cycle(pwm_duty_cycle),
    .out({uio_out, uo_out})
  );

  
  // List all unused inputs to prevent warnings
  
  wire _unused = &{ena, clk, rst_n, 1'b0, uio_in, ui_in[7:3]};

endmodule